//*********************************//
//        Branch Stack             //
//*********************************//

`define  BR_PR_WRONG    1'b0//branch predict wrong
`define  BR_PR_RIGHT    1'b1//branch predict right
